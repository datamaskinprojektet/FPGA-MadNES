`timescale 1ns / 1ps


module top_test_tb();

    parameter CLK_PERIOD = 10;  // 10 ns == 100 MHz

    logic clk;
    logic reset;
    logic [15:0] EBI_AD;
    logic EBI_ALE;
    logic EBI_RE;
    logic EBI_WE;
    logic [2:0] bank_select;
    logic vga_hsync;
    logic vga_vsync;
    logic [3:0] vga_r;
    logic [3:0] vga_g;
    logic [3:0] vga_b;
    logic [50:0] clk_count;

    int fd;

    display_driver dut_display_driver(
    .clk_100m        (clk),             
    .btn_rst         (!reset),             
    .EBI_AD          (EBI_AD),      
    .EBI_ALE         (EBI_ALE),       
    .EBI_RE          (EBI_RE),      
    .EBI_WE          (EBI_WE),      
    .bank_select     (bank_select),            
    .vga_hsync       (vga_hsync),             
    .vga_vsync       (vga_vsync),             
    .vga_r           (vga_r),       
    .vga_g           (vga_g),       
    .vga_b           (vga_b)       
    );                

    always #(CLK_PERIOD / 2) clk = ~clk;

    always @(posedge clk) begin
        clk_count++;
    end


    task resetModule();

        reset = 0;
        clk = 1;
        EBI_AD = 0;
        EBI_ALE = 1;
        EBI_WE = 1;
        EBI_RE = 1;
        bank_select = 0;
        dut_display_driver.OAM.myram_gen[0].myram.memory = '{default:0};
        dut_display_driver.OAM.myram_gen[1].myram.memory = '{default:0};
        //dut_display_driver.TAM.TAM_RAM = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[0].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[1].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[2].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[3].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[4].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[5].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[6].myram.memory = '{default:0};
        //dut_display_driver.SPRITE.myram_gen[7].myram.memory = '{default:0};
        #1;
        reset = 1;
        clk_count = 0;
        #100;
        reset = 0;
        #3000;
    endtask

    task write_oam_data();
        // Generating OAM

        #79.36;
        bank_select = 0;
        EBI_AD = 0;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000100000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 1;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1100000000001000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;

        #79.36;
        EBI_AD = 2;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 3;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1000000000000000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;

        #79.36;

    endtask

    task write_sprite_data();
        // Generating VRAM SPRITE

        #79.36;
        bank_select = 1;
        EBI_AD = 0;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 1;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 2;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 3;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 4;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 5;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 6;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 7;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 8;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 9;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 10;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 11;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 12;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 13;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 14;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 15;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 16;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 17;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 18;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 19;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 20;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 21;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 22;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 23;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 24;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 25;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 26;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 27;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 28;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 29;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 30;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 31;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 32;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 33;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 34;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 35;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 36;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 37;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 38;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 39;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 40;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 41;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 42;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 43;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 44;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 45;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 46;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 47;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 48;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 49;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 50;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 51;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 52;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 53;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 54;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 55;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 56;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 57;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 58;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 59;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 60;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 61;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 62;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 63;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 64;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 65;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 66;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 67;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 68;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 69;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 70;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 71;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 72;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 73;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 74;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 75;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 76;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 77;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 78;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 79;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 80;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 81;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 82;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 83;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 84;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 85;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 86;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 87;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 88;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 89;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 90;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 91;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 92;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 93;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 94;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 95;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 96;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 97;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 98;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 99;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 100;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 101;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 102;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 103;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 104;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 105;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 106;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 107;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 108;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 109;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 110;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 111;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 112;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 113;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 114;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 115;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 116;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 117;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 118;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 119;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 120;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 121;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 122;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 123;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 124;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 125;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 126;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 127;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
    endtask

    task write_pallet_data();
        // Generating Pallet

        #79.36;
        bank_select = 3;
        EBI_AD = 0;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1111111111111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 1;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 2;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1111111111111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 3;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 4;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1111111111111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 5;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 6;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1000010110000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 7;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000010000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 8;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0011001000110010;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 9;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000110010;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 10;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1100100011001000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 11;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011001000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
    endtask

    always @ (posedge dut_display_driver.clk_pix)
    begin
        if(dut_display_driver.de)
        begin
            fd = $fopen("display_data.txt","a"); //Opening file for write
            $fwrite(fd,"%d,%d,%d \n",vga_r,vga_g,vga_b);
            $fclose(fd);
        end
    end

    initial begin
    resetModule();
    $display("topmodule testing");
    write_oam_data();
    write_sprite_data();
    write_pallet_data();
    #18_000_000; // 18 ms (one frame is 16.7 ms)
    $finish;  
        
    end

endmodule

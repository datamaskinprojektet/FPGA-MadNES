`timescale 1ns / 1ps


module top_test_tb();

    parameter CLK_PERIOD = 10;  // 10 ns == 100 MHz

    logic clk;
    logic reset;
    logic [15:0] EBI_AD;
    logic EBI_ALE;
    logic EBI_RE;
    logic EBI_WE;
    logic [2:0] bank_select;
    logic vga_hsync;
    logic vga_vsync;
    logic [3:0] vga_r;
    logic [3:0] vga_g;
    logic [3:0] vga_b;
    logic [50:0] clk_count;



    display_driver dut_display_driver(
    .clk_100m        (clk),             
    .btn_rst         (!reset),             
    .EBI_AD          (EBI_AD),      
    .EBI_ALE         (EBI_ALE),       
    .EBI_RE          (EBI_RE),      
    .EBI_WE          (EBI_WE),      
    .bank_select     (bank_select),            
    .vga_hsync       (vga_hsync),             
    .vga_vsync       (vga_vsync),             
    .vga_r           (vga_r),       
    .vga_g           (vga_g),       
    .vga_b           (vga_b)       
    );                

    always #(CLK_PERIOD / 2) clk = ~clk;

    always @(posedge clk) begin
        clk_count++;
    end


    task resetModule();

        reset = 0;
        clk = 1;
        EBI_AD = 0;
        EBI_ALE = 1;
        EBI_WE = 1;
        EBI_RE = 1;
        bank_select = 0;
        #1;
        reset = 1;
        clk_count = 0;
        #100;
        reset = 0;
        #3000;
    endtask

    task write_oam_data();
        // Generating OAM

        #79.36;
        bank_select = 0;
        EBI_AD = 0;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000101111011;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 1;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1100000000001000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;

        #79.36;
        EBI_AD = 2;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 3;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1000000000000000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;

        #79.36;
    endtask

    task write_sprite_data();
        // Generating VRAM SPRITE

        #79.36;
        bank_select = 1;
        EBI_AD = 0;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 1;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 2;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 3;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 4;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 5;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 6;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 7;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 8;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 9;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 10;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 11;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 12;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 13;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 14;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 15;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 16;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 17;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 18;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 19;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 20;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 21;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 22;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 23;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 24;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 25;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 26;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 27;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 28;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 29;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 30;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 31;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000000001;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
    endtask

    task write_pallet_data();
        // Generating Pallet

        #79.36;
        bank_select = 3;
        EBI_AD = 0;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1111111111111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 1;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 2;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1111111111111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 3;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 4;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1111111111111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 5;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011111111;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 6;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1000010110000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 7;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000010000101;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 8;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0011001000110010;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 9;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000000110010;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 10;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b1100100011001000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
        EBI_AD = 11;
        #1;
        EBI_ALE = 0;
        #1;
        EBI_ALE = 1;
        #1;
        EBI_AD = 16'b0000000011001000;
        #1;
        EBI_WE = 0;
        #1;
        EBI_WE = 1;
        #1;
        #79.36;
    endtask

    initial begin
    resetModule();
    $display("topmodule testing");
    write_oam_data();
    write_sprite_data();
    write_pallet_data();
    #18_000_000; // 18 ms (one frame is 16.7 ms)
    $finish;  
        
    end

endmodule
